package arrint is
	type int_std is array (7 downto 0) of integer;	
end arrint;