package complex is
	type arr2d is array (1 downto 0) of integer;	
end complex;

