library IEEE; 
use IEEE.std_logic_1164.all;

package arr is
	type arr2d is array (2 downto 0,2 downto 0) of std_logic_vector(3 downto 0);
end arr;